../../vhdl-jtag/jtagger.vhd